.title Libre Solar DC/DC converter simulation (without control)

.include "solar/solar_panel_60s.sub"
.include 2n7002k.mod

.model 1N4148 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)
.model MBRS360 D(Is=22.6u Rs=.042 N=1.094 Cjo=480p M=.61 Eg=.69 Xti=2)

* Solar panel
Xpvmodule hs gnd SolarPanel60s Isc=5

* Input filter (high voltage side)
Cin cin gnd 470u
Resr_in cin hs 50m

* Load resistor for testing
*Rload_hs hs gnd 50R

* High-side MOSFET
*D1 sw hs 1N4148
XQhs hs gate_hs sw 2n7002k
Vpwm_hs pwm_hs sw 0 PULSE(0 10 3.2u 10n 10n 6.6u 10u)
Rg_hs gate_hs pwm_hs 10R

* Low-side MOSFET
* MOSFETs pins: D G S S
*M1 bat gate gnd gnd Si7336ADP
*XQ1 0  gate bat 0 MOSFETs_IRFZ44N
XQls sw gate_ls gnd 2n7002k
Vpwm_ls pwm_ls gnd 0 PULSE(0 10 0 10n 10n 3u 10u)
Rg_ls gate_ls pwm_ls 10R

* Main inductor and current measurement shunt
L1 sw shunt 22u
Rshunt shunt bat 2m

* Output filter
Cout cout gnd 220u
Resr_out cout bat 30m

* Battery
Vbat ocvbat gnd dc 12V
Rs_bat ocvbat bat 50m

.control
.options savecurrents
tran 100u 1m
rusage trantime traniter
plot hs sw bat @Rshunt[i]
*destroy all
.endc

.end
