.title Libre Solar DC/DC converter simulation

.include "solar/solar_panel_60s.sub"
.include "adc/ad12.mod"
.include "pwm/pwm.mod"

.model 1N4148 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)
.model MBRS360 D(Is=22.6u Rs=.042 N=1.094 Cjo=480p M=.61 Eg=.69 Xti=2)

* from LTspice
.model Si7336ADP VDMOS(Rg=3.5 Rd=1.2m Rs=800u mtriode=1.9 lambda=0.01 Vto=2.9 Ksubthres=100m Kp=280 Cgdmax=1.6n Cgdmin=200p A=1.5 Cgs=5.2n Cjo=3n M=.5 Is=5p Rb=3m Vds=30 Ron=2.4m Qg=36n)

.model a2d adc_bridge(in_low=0.5 in_high=0.5)
.model d2a dac_bridge

* Interface to Firmware with optional parameters Kp and Ki
.model firmware d_process (process_file="dcdc_utest" process_params=["Kp=10", "Ki=2"])
Acontrol [d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 d10 d11]
+ adclk drst [w0 w1 w2 w3 w4 w5 w6 w7 w8 w9 w10 w11 w12 w13 w14 w15] firmware

* Generate ADC clock
Vadclk aadclk gnd 0 PULSE(0 1 0 1n 1n 156.25n 312.5n)
Aadclk [aadclk] [adclk] a2d

* Generate PWM clock (200 * switching frequency)
Vpwmclk apwmclk gnd 0 PULSE(0 1 0 1n 1n 25n 50n)
Apwmclk [apwmclk] [pwmclk] a2d

* Internal VDD and reference voltage for ADC
Vin vddio 0 DC(3.3)
Vref ref 0 DC(2.048)

* vadc = ADC input (must be below ref)
*Vsolar hs 0 DC(60)
R1 hs vadc 100k
R2 vadc 0 2.2k

* Convert analog reading to digital ADC value
Xad vadc ref vddio adclk d11 d10 d9 d8 d7 d6 d5 d4 d3 d2 d1 d0 ad12

* Generate digital HS and LS PWM signals from compare register value received from control function
Xpwm pwmclk drst w0 w1 w2 w3 w4 w5 w6 w7 w8 w9 w10 w11 w12 w13 w14 w15 dpwm_hs dpwm_ls PWM

* Generate 10V analog PWM signal at high-side gate
Adbridge [dpwm_hs] [pwma_hs] d2a
Bpwmhs pwm_hs sw V=v(pwma_hs)*10

* Generate 10V analog PWM signal at low-side gate
Adbridge2 [dpwm_ls] [pwma_ls] d2a
Bpwmls pwm_ls 0 V=v(pwma_ls)*10

* Solar panel
Xpvmodule hs gnd SolarPanel60s Isc=5

* Input filter (high voltage side)
Cin cin gnd 470u
Resr_in cin hs 50m

* Load resistor for testing
*Rload_hs hs gnd 50R

* High-side MOSFET
Mhs hs gate_hs sw Si7336ADP
Rg_hs gate_hs pwm_hs 20R

* Low-side MOSFET
Mls sw gate_ls gnd Si7336ADP
Rg_ls gate_ls pwm_ls 20R

* Main inductor and current measurement shunt
L1 sw shunt 22u
Rshunt shunt bat 2m

* Output filter
Cout cout gnd 220u
Resr_out cout bat 30m

* Battery
Vbat ocvbat gnd dc 12V
Rs_bat ocvbat bat 50m

.control
.options savecurrents
tran 100u 10m
rusage trantime traniter
plot hs sw bat @Rshunt[i] pwm_ls pwm_hs
*destroy all
.endc

.end
